
`include "apb_if.svh"
`include "uvm_macros.svh"

package prj_pkg;
    import uvm_pkg::*;
    `include "apb_seq_item.svh"
    `include "apb_monitor.svh"
    `include "apb_scoreboard.svh"
    `include "apb_driver.svh"
    `include "apb_sequence.svh"
    `include "apb_sequencer.svh"
    `include "apb_agent.svh"
    `include "apb_env.svh"
    `include "apb_test.svh"
endpackage
